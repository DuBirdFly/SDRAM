// sdr-define
`include "sdr_define.svh"

// sdr-base
`include "IfSdr.sv"
`include "TrSdr.sv"

// sdr-agent
`include "SdrMstrSqr.sv"
`include "SdrMstrChn.sv"
`include "SdrMstrAgt.sv"

// sdr-env
`include "SdrMstrEnv.sv"

// sdr-seq
`include "SdrMstrSeq.sv"
