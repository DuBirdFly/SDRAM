`define VIP_SDR_ADDR_WIDTH  13
`define VIP_SDR_BA_WIDTH     2
`define VIP_SDR_DQ_WIDTH    16
`define VIP_SDR_DM_WIDTH    (`VIP_SDR_DQ_WIDTH / 8)
