typedef uvm_sequencer #(TrSdr) SdrMstrSqr;
