`define VIP_SDR_BA_WIDTH     2

`define VIP_SDR_ADDR_WIDTH  13
`define VIP_SDR_ROW_WIDTH   13
`define VIP_SDR_COL_WIDTH    9

`define VIP_SDR_DQ_WIDTH    16
`define VIP_SDR_DM_WIDTH    (`VIP_SDR_DQ_WIDTH / 8)

`define VIP_SDR_CL_WIDTH     3
`define VIP_SDR_BT_WIDTH     1
`define VIP_SDR_BL_WIDTH     3

// 每一个地址对应 `VIP_SDR_DQ_WIDTH 的数据
`define VIP_NATIVE_ADDR_WIDTH (`VIP_SDR_BA_WIDTH + `VIP_SDR_ROW_WIDTH + `VIP_SDR_COL_WIDTH)
`define VIP_SDR_COL_BASE_ADDR 0
`define VIP_SDR_ROW_BASE_ADDR `VIP_SDR_COL_WIDTH
`define VIP_SDR_BA_BASE_ADDR  (`VIP_SDR_ROW_BASE_ADDR + `VIP_SDR_ROW_WIDTH)
